module sram(cs,oe,we,addr,din,dout);
  input cs;
  input oe;
  input we;
  input [31:0] addr;
  input [31:0] din;
  output reg [31:0] dout;
  
endmodule
